module cpu(

    input wire [31:0] in,
    output reg [31:0] address,
    output reg [31:0] out,
    output reg        we

);

endmodule
